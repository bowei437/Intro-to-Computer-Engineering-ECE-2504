library verilog;
use verilog.vl_types.all;
entity adder4bit_vlg_vec_tst is
end adder4bit_vlg_vec_tst;
