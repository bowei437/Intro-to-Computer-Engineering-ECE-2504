library verilog;
use verilog.vl_types.all;
entity adder1bit_vlg_vec_tst is
end adder1bit_vlg_vec_tst;
