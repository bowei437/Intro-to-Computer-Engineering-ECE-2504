library verilog;
use verilog.vl_types.all;
entity HW3P2_vlg_vec_tst is
end HW3P2_vlg_vec_tst;
