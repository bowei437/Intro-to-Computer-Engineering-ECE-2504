library verilog;
use verilog.vl_types.all;
entity DP3_Spring2015_vlg_vec_tst is
end DP3_Spring2015_vlg_vec_tst;
