library verilog;
use verilog.vl_types.all;
entity DP3_Spring2015_vlg_check_tst is
    port(
        LED             : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end DP3_Spring2015_vlg_check_tst;
