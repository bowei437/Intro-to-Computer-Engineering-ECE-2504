library verilog;
use verilog.vl_types.all;
entity HW41_vlg_check_tst is
    port(
        F1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end HW41_vlg_check_tst;
