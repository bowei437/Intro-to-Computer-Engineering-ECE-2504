library verilog;
use verilog.vl_types.all;
entity DP2_Spring2015_vlg_vec_tst is
end DP2_Spring2015_vlg_vec_tst;
