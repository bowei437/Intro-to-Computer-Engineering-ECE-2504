library verilog;
use verilog.vl_types.all;
entity HW41_vlg_vec_tst is
end HW41_vlg_vec_tst;
