library verilog;
use verilog.vl_types.all;
entity HW3P3 is
    port(
        F1              : out    vl_logic;
        B               : in     vl_logic;
        A               : in     vl_logic;
        D               : in     vl_logic;
        C               : in     vl_logic;
        F2              : out    vl_logic
    );
end HW3P3;
