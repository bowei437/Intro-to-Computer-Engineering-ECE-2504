library verilog;
use verilog.vl_types.all;
entity DP4_ECE2504_vlg_vec_tst is
end DP4_ECE2504_vlg_vec_tst;
