library verilog;
use verilog.vl_types.all;
entity basicmoduleP1_vlg_vec_tst is
end basicmoduleP1_vlg_vec_tst;
