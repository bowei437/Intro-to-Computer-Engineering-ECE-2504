library verilog;
use verilog.vl_types.all;
entity HW3P4_vlg_vec_tst is
end HW3P4_vlg_vec_tst;
